��Q0      �sklearn.ensemble._forest��RandomForestClassifier���)��}�(�base_estimator��sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �_sklearn_version��1.0.2�ub�n_estimators�K
�estimator_params�(hhhhhhhhhht��	bootstrap���	oob_score���n_jobs�NhK*�verbose�K �
warm_start��hN�max_samples�NhhhKhKhKhG        h�auto�hNhG        hG        �feature_names_in_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h)�dtype����O8�����R�(K�|�NNNJ����J����K?t�b�]�(�objawy��wiek��choroby_wsp��wzrost��leki�et�b�n_features_in_�K�
n_outputs_�K�classes_�h(h+K ��h-��R�(KK��h2�i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�
n_classes_�K�base_estimator_�h	�estimators_�]�(h)��}�(hhhhhKhKhKhG        hh$hNhJf��_hG        hNhG        h?Kh@KhAh(h+K ��h-��R�(KK��h2�f8�����R�(KhINNNJ����J����K t�b�C              �?�t�bhMh&�scalar���hHC       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���Kh(h+K ��h-��R�(KK��hH�C       �t�bK��R�}�(hK�
node_count�K	�nodes�h(h+K ��h-��R�(KK	��h2�V56�����R�(Kh6N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hyhHK ��hzhHK��h{hHK��h|hYK��h}hYK ��h~hHK(��hhYK0��uK8KKt�b�B�                              �?�q���?             H@������������������������       �                     (@                           @<ݚ)�?             B@                            @      �?	             (@������������������������       ��eP*L��?             &@������������������������       �                     �?                            @�q�q�?             8@������������������������       ��E��ӭ�?             2@������������������������       �                     @�t�b�values�h(h+K ��h-��R�(KK	KK��hY�C�      7@      9@      (@              &@      9@      @      @      @      @              �?      @      3@      @      *@              @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ�=�KhG        hNhG        h?Kh@KhAh(h+K ��h-��R�(KK��hY�C              �?�t�bhMh^hHC       ���R�hbKhchfKh(h+K ��h-��R�(KK��hH�C       �t�bK��R�}�(hKhpKhqh(h+K ��h-��R�(KK��hx�Bh                           �%g@     ��?             H@                           e@�E��ӭ�?
             2@                          �d@      �?              @������������������������       �                     �?������������������������       �����X�?             @������������������������       �                     $@       
                     @������?             >@       	                   �h@���Q��?             4@������������������������       �      �?             0@������������������������       �                     @������������������������       �                     $@�t�bh�h(h+K ��h-��R�(KKKK��hY�C�      5@      ;@      *@      @      @      @      �?               @      @      $@               @      6@       @      (@       @       @              @              $@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ\bshG        hNhG        h?Kh@KhAh(h+K ��h-��R�(KK��hY�C              �?�t�bhMh^hHC       ���R�hbKhchfKh(h+K ��h-��R�(KK��hH�C       �t�bK��R�}�(hKhpKhqh(h+K ��h-��R�(KK��hx�Bh                            �g@�q���?!             H@                          �E@¦	^_�?             ?@                            @X�Cc�?
             ,@������������������������       �      �?             $@������������������������       �                     @������������������������       �                     1@       
                     @@�0�!��?             1@       	                    @���!pc�?             &@������������������������       �                      @������������������������       ��q�q�?             "@������������������������       �                     @�t�bh�h(h+K ��h-��R�(KKKK��hY�C�      9@      7@      6@      "@      @      "@      @      @              @      1@              @      ,@      @       @               @      @      @              @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ��.hG        hNhG        h?Kh@KhAh(h+K ��h-��R�(KK��hY�C              �?�t�bhMh^hHC       ���R�hbKhchfKh(h+K ��h-��R�(KK��hH�C       �t�bK��R�}�(hKhpKhqh(h+K ��h-��R�(KK��hx�Bh                            �E@r�q��?!             H@                          �0@"pc�
�?             6@������������������������       �                      @                          `h@ףp=
�?             4@������������������������       �"pc�
�?
             &@������������������������       �                     "@       
                    N@8�Z$���?             :@       	                   g@������?
             .@������������������������       �                     $@������������������������       �z�G�z�?             @������������������������       �                     &@�t�bh�h(h+K ��h-��R�(KKKK��hY�C�      :@      6@      @      2@       @               @      2@       @      "@              "@      6@      @      &@      @      $@              �?      @      &@        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJj�c;hG        hNhG        h?Kh@KhAh(h+K ��h-��R�(KK��hY�C              �?�t�bhMh^hHC       ���R�hbKhchfKh(h+K ��h-��R�(KK��hH�C       �t�bK��R�}�(hKhpKhqh(h+K ��h-��R�(KK��hx�B�                            pg@     ��?             H@                          �E@V�a�� �?             =@                            @X�<ݚ�?             "@������������������������       �և���X�?             @������������������������       �                      @                           @P���Q�?             4@������������������������       �        	             1@������������������������       ��q�q�?             @	       
                    7@���y4F�?             3@������������������������       ��q�q�?             @                           N@      �?	             0@������������������������       �$�q-�?             *@������������������������       ��q�q�?             @�t�bh�h(h+K ��h-��R�(KKKK��hY�C�      ;@      5@      7@      @      @      @      @      @               @      3@      �?      1@               @      �?      @      .@       @      �?       @      ,@      �?      (@      �?       @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJGԙGhG        hNhG        h?Kh@KhAh(h+K ��h-��R�(KK��hY�C              �?�t�bhMh^hHC       ���R�hbKhchfKh(h+K ��h-��R�(KK��hH�C       �t�bK��R�}�(hKhpKhqh(h+K ��h-��R�(KK��hx�Bh                              @�q���?             H@                          �h@�!���?             A@                          �E@r֛w���?             ?@������������������������       �X�<ݚ�?             2@������������������������       �        
             *@������������������������       �                     @       
                   0f@؇���X�?             ,@       	                   �d@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     $@�t�bh�h(h+K ��h-��R�(KKKK��hY�C�      9@      7@      7@      &@      7@       @      $@       @      *@                      @       @      (@       @       @               @       @                      $@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ��AhG        hNhG        h?Kh@KhAh(h+K ��h-��R�(KK��hY�C              �?�t�bhMh^hHC       ���R�hbKhchfKh(h+K ��h-��R�(KK��hH�C       �t�bK��R�}�(hKhpKhqh(h+K ��h-��R�(KK��hx�Bh                            �E@r�q��?!             H@                            @��s����?             5@                           @���Q��?	             $@������������������������       �      �?             @������������������������       �      �?             @������������������������       �                     &@                           �?�+$�jP�?             ;@������������������������       �                     @	       
                   �g@      �?             4@������������������������       �                     .@������������������������       �                     @�t�bh�h(h+K ��h-��R�(KKKK��hY�C�      :@      6@      @      1@      @      @      @      @      �?      @              &@      6@      @      @              .@      @      .@                      @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJ,�hG        hNhG        h?Kh@KhAh(h+K ��h-��R�(KK��hY�C              �?�t�bhMh^hHC       ���R�hbKhchfKh(h+K ��h-��R�(KK��hH�C       �t�bK��R�}�(hKhpKhqh(h+K ��h-��R�(KK��hx�Bh                              @�q�q��?             H@                          �h@*;L]n�?             >@                           @$��m��?             :@������������������������       �                     &@������������������������       ����Q��?             .@������������������������       �                     @       
                   0f@�����H�?             2@       	                    @���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     *@�t�bh�h(h+K ��h-��R�(KKKK��hY�C�      3@      =@      1@      *@      1@      "@      &@              @      "@              @       @      0@       @      @       @                      @              *@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJf��'hG        hNhG        h?Kh@KhAh(h+K ��h-��R�(KK��hY�C              �?�t�bhMh^hHC       ���R�hbKhchfKh(h+K ��h-��R�(KK��hH�C       �t�bK��R�}�(hKhpKhqh(h+K ��h-��R�(KK��hx�B�                            �g@r�qG�?             H@                          �E@z�G�z�?            �A@                          @E@և���X�?             @������������������������       �      �?             @������������������������       �                     @                           @ �Cc}�?             <@������������������������       ����7�?             6@������������������������       ��q�q�?             @	       
                    @�θ�?
             *@������������������������       �                     @                          �;@�q�q�?             "@������������������������       �      �?             @������������������������       �                     @�t�bh�h(h+K ��h-��R�(KKKK��hY�C�      ?@      1@      <@      @      @      @      @      �?              @      9@      @      5@      �?      @       @      @      $@              @      @      @      @      @              @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh$hNhJy"rhG        hNhG        h?Kh@KhAh(h+K ��h-��R�(KK��hY�C              �?�t�bhMh^hHC       ���R�hbKhchfKh(h+K ��h-��R�(KK��hH�C       �t�bK��R�}�(hKhpKhqh(h+K ��h-��R�(KK��hx�Bh                              �?      �?             H@                         y�H@�IєX�?	             1@                           @z�G�z�?             @������������������������       �      �?              @������������������������       �                     @������������������������       �                     (@                           '@r֛w���?             ?@������������������������       �                      @	       
                  �%g@V�a�� �?             =@������������������������       ��q�q�?             (@������������������������       ��t����?             1@�t�bh�h(h+K ��h-��R�(KKKK��hY�C�      8@      8@      0@      �?      @      �?      �?      �?      @              (@               @      7@       @              @      7@      @       @       @      .@�t�bubhhubehhub.